module main

struct Food {
	pos			Position
}
